library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 14; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0efc287",
    12 => x"86c0c84e",
    13 => x"49f0efc2",
    14 => x"48fcdcc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f1e2",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34972",
    82 => x"c27c7199",
    83 => x"05bffcdc",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"c329d849",
    88 => x"7c7199ff",
    89 => x"d04966d0",
    90 => x"99ffc329",
    91 => x"66d07c71",
    92 => x"c329c849",
    93 => x"7c7199ff",
    94 => x"c34966d0",
    95 => x"7c7199ff",
    96 => x"29d04972",
    97 => x"7199ffc3",
    98 => x"c94b6c7c",
    99 => x"c34dfff0",
   100 => x"d005abff",
   101 => x"7cffc387",
   102 => x"8dc14b6c",
   103 => x"c387c602",
   104 => x"f002abff",
   105 => x"fe487387",
   106 => x"c01e87c7",
   107 => x"48d4ff49",
   108 => x"c178ffc3",
   109 => x"b7c8c381",
   110 => x"87f104a9",
   111 => x"731e4f26",
   112 => x"c487e71e",
   113 => x"c04bdff8",
   114 => x"f0ffc01e",
   115 => x"fd49f7c1",
   116 => x"86c487e7",
   117 => x"c005a8c1",
   118 => x"d4ff87ea",
   119 => x"78ffc348",
   120 => x"c0c0c0c1",
   121 => x"c01ec0c0",
   122 => x"e9c1f0e1",
   123 => x"87c9fd49",
   124 => x"987086c4",
   125 => x"ff87ca05",
   126 => x"ffc348d4",
   127 => x"cb48c178",
   128 => x"87e6fe87",
   129 => x"fe058bc1",
   130 => x"48c087fd",
   131 => x"1e87e6fc",
   132 => x"d4ff1e73",
   133 => x"78ffc348",
   134 => x"1ec04bd3",
   135 => x"c1f0ffc0",
   136 => x"d4fc49c1",
   137 => x"7086c487",
   138 => x"87ca0598",
   139 => x"c348d4ff",
   140 => x"48c178ff",
   141 => x"f1fd87cb",
   142 => x"058bc187",
   143 => x"c087dbff",
   144 => x"87f1fb48",
   145 => x"5c5b5e0e",
   146 => x"4cd4ff0e",
   147 => x"c687dbfd",
   148 => x"e1c01eea",
   149 => x"49c8c1f0",
   150 => x"c487defb",
   151 => x"02a8c186",
   152 => x"eafe87c8",
   153 => x"c148c087",
   154 => x"dafa87e2",
   155 => x"cf497087",
   156 => x"c699ffff",
   157 => x"c802a9ea",
   158 => x"87d3fe87",
   159 => x"cbc148c0",
   160 => x"7cffc387",
   161 => x"fc4bf1c0",
   162 => x"987087f4",
   163 => x"87ebc002",
   164 => x"ffc01ec0",
   165 => x"49fac1f0",
   166 => x"c487defa",
   167 => x"05987086",
   168 => x"ffc387d9",
   169 => x"c3496c7c",
   170 => x"7c7c7cff",
   171 => x"99c0c17c",
   172 => x"c187c402",
   173 => x"c087d548",
   174 => x"c287d148",
   175 => x"87c405ab",
   176 => x"87c848c0",
   177 => x"fe058bc1",
   178 => x"48c087fd",
   179 => x"1e87e4f9",
   180 => x"dcc21e73",
   181 => x"78c148fc",
   182 => x"d0ff4bc7",
   183 => x"fb78c248",
   184 => x"d0ff87c8",
   185 => x"c078c348",
   186 => x"d0e5c01e",
   187 => x"f949c0c1",
   188 => x"86c487c7",
   189 => x"c105a8c1",
   190 => x"abc24b87",
   191 => x"c087c505",
   192 => x"87f9c048",
   193 => x"ff058bc1",
   194 => x"f7fc87d0",
   195 => x"c0ddc287",
   196 => x"05987058",
   197 => x"1ec187cd",
   198 => x"c1f0ffc0",
   199 => x"d8f849d0",
   200 => x"ff86c487",
   201 => x"ffc348d4",
   202 => x"87dec478",
   203 => x"58c4ddc2",
   204 => x"c248d0ff",
   205 => x"48d4ff78",
   206 => x"c178ffc3",
   207 => x"87f5f748",
   208 => x"5c5b5e0e",
   209 => x"4a710e5d",
   210 => x"ff4dffc3",
   211 => x"7c754cd4",
   212 => x"c448d0ff",
   213 => x"7c7578c3",
   214 => x"ffc01e72",
   215 => x"49d8c1f0",
   216 => x"c487d6f7",
   217 => x"02987086",
   218 => x"48c187c5",
   219 => x"7587f0c0",
   220 => x"7cfec37c",
   221 => x"d41ec0c8",
   222 => x"faf44966",
   223 => x"7586c487",
   224 => x"757c757c",
   225 => x"e0dad87c",
   226 => x"6c7c754b",
   227 => x"c5059949",
   228 => x"058bc187",
   229 => x"7c7587f3",
   230 => x"c248d0ff",
   231 => x"f648c078",
   232 => x"5e0e87cf",
   233 => x"0e5d5c5b",
   234 => x"4cc04b71",
   235 => x"dfcdeec5",
   236 => x"48d4ff4a",
   237 => x"6878ffc3",
   238 => x"a9fec349",
   239 => x"87fdc005",
   240 => x"9b734d70",
   241 => x"d087cc02",
   242 => x"49731e66",
   243 => x"c487cff4",
   244 => x"ff87d686",
   245 => x"d1c448d0",
   246 => x"7dffc378",
   247 => x"c14866d0",
   248 => x"58a6d488",
   249 => x"f0059870",
   250 => x"48d4ff87",
   251 => x"7878ffc3",
   252 => x"c5059b73",
   253 => x"48d0ff87",
   254 => x"4ac178d0",
   255 => x"058ac14c",
   256 => x"7487eefe",
   257 => x"87e9f448",
   258 => x"711e731e",
   259 => x"ff4bc04a",
   260 => x"ffc348d4",
   261 => x"48d0ff78",
   262 => x"ff78c3c4",
   263 => x"ffc348d4",
   264 => x"c01e7278",
   265 => x"d1c1f0ff",
   266 => x"87cdf449",
   267 => x"987086c4",
   268 => x"c887d205",
   269 => x"66cc1ec0",
   270 => x"87e6fd49",
   271 => x"4b7086c4",
   272 => x"c248d0ff",
   273 => x"f3487378",
   274 => x"5e0e87eb",
   275 => x"0e5d5c5b",
   276 => x"ffc01ec0",
   277 => x"49c9c1f0",
   278 => x"d287def3",
   279 => x"c4ddc21e",
   280 => x"87fefc49",
   281 => x"4cc086c8",
   282 => x"b7d284c1",
   283 => x"87f804ac",
   284 => x"97c4ddc2",
   285 => x"c0c349bf",
   286 => x"a9c0c199",
   287 => x"87e7c005",
   288 => x"97cbddc2",
   289 => x"31d049bf",
   290 => x"97ccddc2",
   291 => x"32c84abf",
   292 => x"ddc2b172",
   293 => x"4abf97cd",
   294 => x"cf4c71b1",
   295 => x"9cffffff",
   296 => x"34ca84c1",
   297 => x"c287e7c1",
   298 => x"bf97cddd",
   299 => x"c631c149",
   300 => x"ceddc299",
   301 => x"c74abf97",
   302 => x"b1722ab7",
   303 => x"97c9ddc2",
   304 => x"cf4d4abf",
   305 => x"caddc29d",
   306 => x"c34abf97",
   307 => x"c232ca9a",
   308 => x"bf97cbdd",
   309 => x"7333c24b",
   310 => x"ccddc2b2",
   311 => x"c34bbf97",
   312 => x"b7c69bc0",
   313 => x"c2b2732b",
   314 => x"7148c181",
   315 => x"c1497030",
   316 => x"70307548",
   317 => x"c14c724d",
   318 => x"c8947184",
   319 => x"06adb7c0",
   320 => x"34c187cc",
   321 => x"c0c82db7",
   322 => x"ff01adb7",
   323 => x"487487f4",
   324 => x"0e87def0",
   325 => x"5d5c5b5e",
   326 => x"c286f80e",
   327 => x"c048eae5",
   328 => x"e2ddc278",
   329 => x"fb49c01e",
   330 => x"86c487de",
   331 => x"c5059870",
   332 => x"c948c087",
   333 => x"4dc087ce",
   334 => x"f2c07ec1",
   335 => x"c249bfec",
   336 => x"714ad8de",
   337 => x"e0ec4bc8",
   338 => x"05987087",
   339 => x"7ec087c2",
   340 => x"bfe8f2c0",
   341 => x"f4dec249",
   342 => x"4bc8714a",
   343 => x"7087caec",
   344 => x"87c20598",
   345 => x"026e7ec0",
   346 => x"c287fdc0",
   347 => x"4dbfe8e4",
   348 => x"9fe0e5c2",
   349 => x"c5487ebf",
   350 => x"05a8ead6",
   351 => x"e4c287c7",
   352 => x"ce4dbfe8",
   353 => x"ca486e87",
   354 => x"02a8d5e9",
   355 => x"48c087c5",
   356 => x"c287f1c7",
   357 => x"751ee2dd",
   358 => x"87ecf949",
   359 => x"987086c4",
   360 => x"c087c505",
   361 => x"87dcc748",
   362 => x"bfe8f2c0",
   363 => x"f4dec249",
   364 => x"4bc8714a",
   365 => x"7087f2ea",
   366 => x"87c80598",
   367 => x"48eae5c2",
   368 => x"87da78c1",
   369 => x"bfecf2c0",
   370 => x"d8dec249",
   371 => x"4bc8714a",
   372 => x"7087d6ea",
   373 => x"c5c00298",
   374 => x"c648c087",
   375 => x"e5c287e6",
   376 => x"49bf97e0",
   377 => x"05a9d5c1",
   378 => x"c287cdc0",
   379 => x"bf97e1e5",
   380 => x"a9eac249",
   381 => x"87c5c002",
   382 => x"c7c648c0",
   383 => x"e2ddc287",
   384 => x"487ebf97",
   385 => x"02a8e9c3",
   386 => x"6e87cec0",
   387 => x"a8ebc348",
   388 => x"87c5c002",
   389 => x"ebc548c0",
   390 => x"edddc287",
   391 => x"9949bf97",
   392 => x"87ccc005",
   393 => x"97eeddc2",
   394 => x"a9c249bf",
   395 => x"87c5c002",
   396 => x"cfc548c0",
   397 => x"efddc287",
   398 => x"c248bf97",
   399 => x"7058e6e5",
   400 => x"88c1484c",
   401 => x"58eae5c2",
   402 => x"97f0ddc2",
   403 => x"817549bf",
   404 => x"97f1ddc2",
   405 => x"32c84abf",
   406 => x"c27ea172",
   407 => x"6e48f7e9",
   408 => x"f2ddc278",
   409 => x"c848bf97",
   410 => x"e5c258a6",
   411 => x"c202bfea",
   412 => x"f2c087d4",
   413 => x"c249bfe8",
   414 => x"714af4de",
   415 => x"e8e74bc8",
   416 => x"02987087",
   417 => x"c087c5c0",
   418 => x"87f8c348",
   419 => x"bfe2e5c2",
   420 => x"cbeac24c",
   421 => x"c7dec25c",
   422 => x"c849bf97",
   423 => x"c6dec231",
   424 => x"a14abf97",
   425 => x"c8dec249",
   426 => x"d04abf97",
   427 => x"49a17232",
   428 => x"97c9dec2",
   429 => x"32d84abf",
   430 => x"c449a172",
   431 => x"e9c29166",
   432 => x"c281bff7",
   433 => x"c259ffe9",
   434 => x"bf97cfde",
   435 => x"c232c84a",
   436 => x"bf97cede",
   437 => x"c24aa24b",
   438 => x"bf97d0de",
   439 => x"7333d04b",
   440 => x"dec24aa2",
   441 => x"4bbf97d1",
   442 => x"33d89bcf",
   443 => x"c24aa273",
   444 => x"c25ac3ea",
   445 => x"4abfffe9",
   446 => x"92748ac2",
   447 => x"48c3eac2",
   448 => x"c178a172",
   449 => x"ddc287ca",
   450 => x"49bf97f4",
   451 => x"ddc231c8",
   452 => x"4abf97f3",
   453 => x"e5c249a1",
   454 => x"e5c259f2",
   455 => x"c549bfee",
   456 => x"81ffc731",
   457 => x"eac229c9",
   458 => x"ddc259cb",
   459 => x"4abf97f9",
   460 => x"ddc232c8",
   461 => x"4bbf97f8",
   462 => x"66c44aa2",
   463 => x"c2826e92",
   464 => x"c25ac7ea",
   465 => x"c048ffe9",
   466 => x"fbe9c278",
   467 => x"78a17248",
   468 => x"48cbeac2",
   469 => x"bfffe9c2",
   470 => x"cfeac278",
   471 => x"c3eac248",
   472 => x"e5c278bf",
   473 => x"c002bfea",
   474 => x"487487c9",
   475 => x"7e7030c4",
   476 => x"c287c9c0",
   477 => x"48bfc7ea",
   478 => x"7e7030c4",
   479 => x"48eee5c2",
   480 => x"48c1786e",
   481 => x"4d268ef8",
   482 => x"4b264c26",
   483 => x"5e0e4f26",
   484 => x"0e5d5c5b",
   485 => x"e5c24a71",
   486 => x"cb02bfea",
   487 => x"c74b7287",
   488 => x"c14c722b",
   489 => x"87c99cff",
   490 => x"2bc84b72",
   491 => x"ffc34c72",
   492 => x"f7e9c29c",
   493 => x"f2c083bf",
   494 => x"02abbfe4",
   495 => x"f2c087d9",
   496 => x"ddc25be8",
   497 => x"49731ee2",
   498 => x"c487fdf0",
   499 => x"05987086",
   500 => x"48c087c5",
   501 => x"c287e6c0",
   502 => x"02bfeae5",
   503 => x"497487d2",
   504 => x"ddc291c4",
   505 => x"4d6981e2",
   506 => x"ffffffcf",
   507 => x"87cb9dff",
   508 => x"91c24974",
   509 => x"81e2ddc2",
   510 => x"754d699f",
   511 => x"87c6fe48",
   512 => x"5c5b5e0e",
   513 => x"86f80e5d",
   514 => x"059c4c71",
   515 => x"48c087c5",
   516 => x"c887c1c3",
   517 => x"c0487ea4",
   518 => x"0266d878",
   519 => x"66d887c7",
   520 => x"c505bf97",
   521 => x"c248c087",
   522 => x"1ec087ea",
   523 => x"ca4949c1",
   524 => x"86c487d7",
   525 => x"029d4d70",
   526 => x"c287c2c1",
   527 => x"d84af2e5",
   528 => x"c9e04966",
   529 => x"02987087",
   530 => x"7587f2c0",
   531 => x"4966d84a",
   532 => x"eee04bcb",
   533 => x"02987087",
   534 => x"c087e2c0",
   535 => x"029d751e",
   536 => x"a6c887c7",
   537 => x"c578c048",
   538 => x"48a6c887",
   539 => x"66c878c1",
   540 => x"87d5c949",
   541 => x"4d7086c4",
   542 => x"fefe059d",
   543 => x"029d7587",
   544 => x"dc87cfc1",
   545 => x"486e49a5",
   546 => x"a5da7869",
   547 => x"48a6c449",
   548 => x"9f78a4c4",
   549 => x"66c44869",
   550 => x"e5c27808",
   551 => x"d202bfea",
   552 => x"49a5d487",
   553 => x"c049699f",
   554 => x"7199ffff",
   555 => x"7030d048",
   556 => x"c087c27e",
   557 => x"48496e7e",
   558 => x"80bf66c4",
   559 => x"780866c4",
   560 => x"a4cc7cc0",
   561 => x"bf66c449",
   562 => x"49a4d079",
   563 => x"48c179c0",
   564 => x"48c087c2",
   565 => x"edfa8ef8",
   566 => x"5b5e0e87",
   567 => x"710e5d5c",
   568 => x"c1029c4c",
   569 => x"a4c887ca",
   570 => x"c1026949",
   571 => x"66d087c2",
   572 => x"82496c4a",
   573 => x"d05aa6d4",
   574 => x"c2b94d66",
   575 => x"4abfe6e5",
   576 => x"9972baff",
   577 => x"c0029971",
   578 => x"a4c487e4",
   579 => x"f9496b4b",
   580 => x"7b7087fc",
   581 => x"bfe2e5c2",
   582 => x"71816c49",
   583 => x"c2b9757c",
   584 => x"4abfe6e5",
   585 => x"9972baff",
   586 => x"ff059971",
   587 => x"7c7587dc",
   588 => x"1e87d3f9",
   589 => x"4b711e73",
   590 => x"87c7029b",
   591 => x"6949a3c8",
   592 => x"c087c505",
   593 => x"87f7c048",
   594 => x"bffbe9c2",
   595 => x"49a3c44a",
   596 => x"89c24969",
   597 => x"bfe2e5c2",
   598 => x"4aa27191",
   599 => x"bfe6e5c2",
   600 => x"71996b49",
   601 => x"f2c04aa2",
   602 => x"66c85ae8",
   603 => x"ea49721e",
   604 => x"86c487d6",
   605 => x"c4059870",
   606 => x"c248c087",
   607 => x"f848c187",
   608 => x"731e87c8",
   609 => x"9b4b711e",
   610 => x"c887c702",
   611 => x"056949a3",
   612 => x"48c087c5",
   613 => x"c287f7c0",
   614 => x"4abffbe9",
   615 => x"6949a3c4",
   616 => x"c289c249",
   617 => x"91bfe2e5",
   618 => x"c24aa271",
   619 => x"49bfe6e5",
   620 => x"a271996b",
   621 => x"e8f2c04a",
   622 => x"1e66c85a",
   623 => x"ffe54972",
   624 => x"7086c487",
   625 => x"87c40598",
   626 => x"87c248c0",
   627 => x"f9f648c1",
   628 => x"5b5e0e87",
   629 => x"1e0e5d5c",
   630 => x"66d44b71",
   631 => x"029b734d",
   632 => x"c887ccc1",
   633 => x"026949a3",
   634 => x"d087c4c1",
   635 => x"e5c24ca3",
   636 => x"ff49bfe6",
   637 => x"994a6cb9",
   638 => x"a966d47e",
   639 => x"c087cd06",
   640 => x"a3cc7c7b",
   641 => x"49a3c44a",
   642 => x"87ca796a",
   643 => x"c0f84972",
   644 => x"4d66d499",
   645 => x"49758d71",
   646 => x"1e7129c9",
   647 => x"f8fa4973",
   648 => x"e2ddc287",
   649 => x"fc49731e",
   650 => x"86c887c9",
   651 => x"267c66d4",
   652 => x"1e87d3f5",
   653 => x"4b711e73",
   654 => x"e4c0029b",
   655 => x"cfeac287",
   656 => x"c24a735b",
   657 => x"e2e5c28a",
   658 => x"c29249bf",
   659 => x"48bffbe9",
   660 => x"eac28072",
   661 => x"487158d3",
   662 => x"e5c230c4",
   663 => x"edc058f2",
   664 => x"cbeac287",
   665 => x"ffe9c248",
   666 => x"eac278bf",
   667 => x"eac248cf",
   668 => x"c278bfc3",
   669 => x"02bfeae5",
   670 => x"e5c287c9",
   671 => x"c449bfe2",
   672 => x"c287c731",
   673 => x"49bfc7ea",
   674 => x"e5c231c4",
   675 => x"f9f359f2",
   676 => x"5b5e0e87",
   677 => x"4a710e5c",
   678 => x"9a724bc0",
   679 => x"87e1c002",
   680 => x"9f49a2da",
   681 => x"e5c24b69",
   682 => x"cf02bfea",
   683 => x"49a2d487",
   684 => x"4c49699f",
   685 => x"9cffffc0",
   686 => x"87c234d0",
   687 => x"49744cc0",
   688 => x"fd4973b3",
   689 => x"fff287ed",
   690 => x"5b5e0e87",
   691 => x"f40e5d5c",
   692 => x"c04a7186",
   693 => x"029a727e",
   694 => x"ddc287d8",
   695 => x"78c048de",
   696 => x"48d6ddc2",
   697 => x"bfcfeac2",
   698 => x"daddc278",
   699 => x"cbeac248",
   700 => x"e5c278bf",
   701 => x"50c048ff",
   702 => x"bfeee5c2",
   703 => x"deddc249",
   704 => x"aa714abf",
   705 => x"87c9c403",
   706 => x"99cf4972",
   707 => x"87e9c005",
   708 => x"48e4f2c0",
   709 => x"bfd6ddc2",
   710 => x"e2ddc278",
   711 => x"d6ddc21e",
   712 => x"ddc249bf",
   713 => x"a1c148d6",
   714 => x"dbe37178",
   715 => x"c086c487",
   716 => x"c248e0f2",
   717 => x"cc78e2dd",
   718 => x"e0f2c087",
   719 => x"e0c048bf",
   720 => x"e4f2c080",
   721 => x"deddc258",
   722 => x"80c148bf",
   723 => x"58e2ddc2",
   724 => x"000ca027",
   725 => x"bf97bf00",
   726 => x"c2029d4d",
   727 => x"e5c387e3",
   728 => x"dcc202ad",
   729 => x"e0f2c087",
   730 => x"a3cb4bbf",
   731 => x"cf4c1149",
   732 => x"d2c105ac",
   733 => x"df497587",
   734 => x"cd89c199",
   735 => x"f2e5c291",
   736 => x"4aa3c181",
   737 => x"a3c35112",
   738 => x"c551124a",
   739 => x"51124aa3",
   740 => x"124aa3c7",
   741 => x"4aa3c951",
   742 => x"a3ce5112",
   743 => x"d051124a",
   744 => x"51124aa3",
   745 => x"124aa3d2",
   746 => x"4aa3d451",
   747 => x"a3d65112",
   748 => x"d851124a",
   749 => x"51124aa3",
   750 => x"124aa3dc",
   751 => x"4aa3de51",
   752 => x"7ec15112",
   753 => x"7487fac0",
   754 => x"0599c849",
   755 => x"7487ebc0",
   756 => x"0599d049",
   757 => x"66dc87d1",
   758 => x"87cbc002",
   759 => x"66dc4973",
   760 => x"0298700f",
   761 => x"6e87d3c0",
   762 => x"87c6c005",
   763 => x"48f2e5c2",
   764 => x"f2c050c0",
   765 => x"c248bfe0",
   766 => x"e5c287e1",
   767 => x"50c048ff",
   768 => x"eee5c27e",
   769 => x"ddc249bf",
   770 => x"714abfde",
   771 => x"f7fb04aa",
   772 => x"cfeac287",
   773 => x"c8c005bf",
   774 => x"eae5c287",
   775 => x"f8c102bf",
   776 => x"daddc287",
   777 => x"e5ed49bf",
   778 => x"c2497087",
   779 => x"c459dedd",
   780 => x"ddc248a6",
   781 => x"c278bfda",
   782 => x"02bfeae5",
   783 => x"c487d8c0",
   784 => x"ffcf4966",
   785 => x"99f8ffff",
   786 => x"c5c002a9",
   787 => x"c04cc087",
   788 => x"4cc187e1",
   789 => x"c487dcc0",
   790 => x"ffcf4966",
   791 => x"02a999f8",
   792 => x"c887c8c0",
   793 => x"78c048a6",
   794 => x"c887c5c0",
   795 => x"78c148a6",
   796 => x"744c66c8",
   797 => x"e0c0059c",
   798 => x"4966c487",
   799 => x"e5c289c2",
   800 => x"914abfe2",
   801 => x"bffbe9c2",
   802 => x"d6ddc24a",
   803 => x"78a17248",
   804 => x"48deddc2",
   805 => x"dff978c0",
   806 => x"f448c087",
   807 => x"87e6eb8e",
   808 => x"00000000",
   809 => x"ffffffff",
   810 => x"00000cb0",
   811 => x"00000cb9",
   812 => x"33544146",
   813 => x"20202032",
   814 => x"54414600",
   815 => x"20203631",
   816 => x"ff1e0020",
   817 => x"ffc348d4",
   818 => x"26486878",
   819 => x"d4ff1e4f",
   820 => x"78ffc348",
   821 => x"c048d0ff",
   822 => x"d4ff78e1",
   823 => x"c278d448",
   824 => x"ff48d3ea",
   825 => x"2650bfd4",
   826 => x"d0ff1e4f",
   827 => x"78e0c048",
   828 => x"ff1e4f26",
   829 => x"497087cc",
   830 => x"87c60299",
   831 => x"05a9fbc0",
   832 => x"487187f1",
   833 => x"5e0e4f26",
   834 => x"710e5c5b",
   835 => x"fe4cc04b",
   836 => x"497087f0",
   837 => x"f9c00299",
   838 => x"a9ecc087",
   839 => x"87f2c002",
   840 => x"02a9fbc0",
   841 => x"cc87ebc0",
   842 => x"03acb766",
   843 => x"66d087c7",
   844 => x"7187c202",
   845 => x"02997153",
   846 => x"84c187c2",
   847 => x"7087c3fe",
   848 => x"cd029949",
   849 => x"a9ecc087",
   850 => x"c087c702",
   851 => x"ff05a9fb",
   852 => x"66d087d5",
   853 => x"c087c302",
   854 => x"ecc07b97",
   855 => x"87c405a9",
   856 => x"87c54a74",
   857 => x"0ac04a74",
   858 => x"c248728a",
   859 => x"264d2687",
   860 => x"264b264c",
   861 => x"c9fd1e4f",
   862 => x"4a497087",
   863 => x"04aaf0c0",
   864 => x"f9c087c9",
   865 => x"87c301aa",
   866 => x"c18af0c0",
   867 => x"c904aac1",
   868 => x"aadac187",
   869 => x"c087c301",
   870 => x"48728af7",
   871 => x"5e0e4f26",
   872 => x"710e5c5b",
   873 => x"4bd4ff4a",
   874 => x"e7c04972",
   875 => x"9c4c7087",
   876 => x"c187c202",
   877 => x"48d0ff8c",
   878 => x"d5c178c5",
   879 => x"c649747b",
   880 => x"d2e4c131",
   881 => x"484abf97",
   882 => x"7b70b071",
   883 => x"c448d0ff",
   884 => x"87dbfe78",
   885 => x"5c5b5e0e",
   886 => x"86f80e5d",
   887 => x"7ec04c71",
   888 => x"c087eafb",
   889 => x"c1fac04b",
   890 => x"c049bf97",
   891 => x"87cf04a9",
   892 => x"c187fffb",
   893 => x"c1fac083",
   894 => x"ab49bf97",
   895 => x"c087f106",
   896 => x"bf97c1fa",
   897 => x"fa87cf02",
   898 => x"497087f8",
   899 => x"87c60299",
   900 => x"05a9ecc0",
   901 => x"4bc087f1",
   902 => x"7087e7fa",
   903 => x"87e2fa4d",
   904 => x"fa58a6c8",
   905 => x"4a7087dc",
   906 => x"a4c883c1",
   907 => x"49699749",
   908 => x"87c702ad",
   909 => x"05adffc0",
   910 => x"c987e7c0",
   911 => x"699749a4",
   912 => x"a966c449",
   913 => x"4887c702",
   914 => x"05a8ffc0",
   915 => x"a4ca87d4",
   916 => x"49699749",
   917 => x"87c602aa",
   918 => x"05aaffc0",
   919 => x"7ec187c4",
   920 => x"ecc087d0",
   921 => x"87c602ad",
   922 => x"05adfbc0",
   923 => x"4bc087c4",
   924 => x"026e7ec1",
   925 => x"f987e1fe",
   926 => x"487387ef",
   927 => x"ecfb8ef8",
   928 => x"5e0e0087",
   929 => x"0e5d5c5b",
   930 => x"4d7186f8",
   931 => x"754bd4ff",
   932 => x"d8eac21e",
   933 => x"87e8e549",
   934 => x"987086c4",
   935 => x"87ccc402",
   936 => x"c148a6c4",
   937 => x"78bfd4e4",
   938 => x"f1fb4975",
   939 => x"48d0ff87",
   940 => x"d6c178c5",
   941 => x"754ac07b",
   942 => x"7b1149a2",
   943 => x"b7cb82c1",
   944 => x"87f304aa",
   945 => x"ffc34acc",
   946 => x"c082c17b",
   947 => x"04aab7e0",
   948 => x"d0ff87f4",
   949 => x"c378c448",
   950 => x"78c57bff",
   951 => x"c17bd3c1",
   952 => x"6678c47b",
   953 => x"a8b7c048",
   954 => x"87f0c206",
   955 => x"bfe0eac2",
   956 => x"4866c44c",
   957 => x"a6c88874",
   958 => x"029c7458",
   959 => x"c287f9c1",
   960 => x"c87ee2dd",
   961 => x"c08c4dc0",
   962 => x"c603acb7",
   963 => x"a4c0c887",
   964 => x"c24cc04d",
   965 => x"bf97d3ea",
   966 => x"0299d049",
   967 => x"1ec087d1",
   968 => x"49d8eac2",
   969 => x"c487cce8",
   970 => x"4a497086",
   971 => x"c287eec0",
   972 => x"c21ee2dd",
   973 => x"e749d8ea",
   974 => x"86c487f9",
   975 => x"ff4a4970",
   976 => x"c5c848d0",
   977 => x"7bd4c178",
   978 => x"7bbf976e",
   979 => x"80c1486e",
   980 => x"8dc17e70",
   981 => x"87f0ff05",
   982 => x"c448d0ff",
   983 => x"059a7278",
   984 => x"48c087c5",
   985 => x"c187c7c1",
   986 => x"d8eac21e",
   987 => x"87e9e549",
   988 => x"9c7486c4",
   989 => x"87c7fe05",
   990 => x"c04866c4",
   991 => x"d106a8b7",
   992 => x"d8eac287",
   993 => x"d078c048",
   994 => x"f478c080",
   995 => x"e4eac280",
   996 => x"66c478bf",
   997 => x"a8b7c048",
   998 => x"87d0fd01",
   999 => x"c548d0ff",
  1000 => x"7bd3c178",
  1001 => x"78c47bc0",
  1002 => x"87c248c1",
  1003 => x"8ef848c0",
  1004 => x"4c264d26",
  1005 => x"4f264b26",
  1006 => x"5c5b5e0e",
  1007 => x"711e0e5d",
  1008 => x"4d4cc04b",
  1009 => x"e8c004ab",
  1010 => x"d4f7c087",
  1011 => x"029d751e",
  1012 => x"4ac087c4",
  1013 => x"4ac187c2",
  1014 => x"eceb4972",
  1015 => x"7086c487",
  1016 => x"6e84c17e",
  1017 => x"7387c205",
  1018 => x"7385c14c",
  1019 => x"d8ff06ac",
  1020 => x"26486e87",
  1021 => x"0e87f9fe",
  1022 => x"0e5c5b5e",
  1023 => x"66cc4b71",
  1024 => x"4c87d802",
  1025 => x"028cf0c0",
  1026 => x"4a7487d8",
  1027 => x"d1028ac1",
  1028 => x"cd028a87",
  1029 => x"c9028a87",
  1030 => x"7387d987",
  1031 => x"87e2f949",
  1032 => x"1e7487d2",
  1033 => x"d8c149c0",
  1034 => x"1e7487ff",
  1035 => x"d8c14973",
  1036 => x"86c887f7",
  1037 => x"0e87fbfd",
  1038 => x"5d5c5b5e",
  1039 => x"4c711e0e",
  1040 => x"c291de49",
  1041 => x"714dc0eb",
  1042 => x"026d9785",
  1043 => x"c287ddc1",
  1044 => x"4abfecea",
  1045 => x"49728274",
  1046 => x"7087ddfd",
  1047 => x"0298487e",
  1048 => x"c287f2c0",
  1049 => x"704bf4ea",
  1050 => x"ff49cb4a",
  1051 => x"7487f8c0",
  1052 => x"c193cb4b",
  1053 => x"c483e6e4",
  1054 => x"f0c2c183",
  1055 => x"c149747b",
  1056 => x"7587ccc1",
  1057 => x"d3e4c17b",
  1058 => x"1e49bf97",
  1059 => x"49f4eac2",
  1060 => x"c487e4fd",
  1061 => x"c1497486",
  1062 => x"c087f4c0",
  1063 => x"d3c2c149",
  1064 => x"d4eac287",
  1065 => x"c178c048",
  1066 => x"87dede49",
  1067 => x"87c0fc26",
  1068 => x"64616f4c",
  1069 => x"2e676e69",
  1070 => x"0e002e2e",
  1071 => x"0e5c5b5e",
  1072 => x"c24a4b71",
  1073 => x"82bfecea",
  1074 => x"ebfb4972",
  1075 => x"9c4c7087",
  1076 => x"4987c402",
  1077 => x"c287fae6",
  1078 => x"c048ecea",
  1079 => x"dd49c178",
  1080 => x"cdfb87e8",
  1081 => x"5b5e0e87",
  1082 => x"f40e5d5c",
  1083 => x"e2ddc286",
  1084 => x"c44cc04d",
  1085 => x"78c048a6",
  1086 => x"bfeceac2",
  1087 => x"06a9c049",
  1088 => x"c287c1c1",
  1089 => x"9848e2dd",
  1090 => x"87f8c002",
  1091 => x"1ed4f7c0",
  1092 => x"c70266c8",
  1093 => x"48a6c487",
  1094 => x"87c578c0",
  1095 => x"c148a6c4",
  1096 => x"4966c478",
  1097 => x"c487e2e6",
  1098 => x"c14d7086",
  1099 => x"4866c484",
  1100 => x"a6c880c1",
  1101 => x"eceac258",
  1102 => x"03ac49bf",
  1103 => x"9d7587c6",
  1104 => x"87c8ff05",
  1105 => x"9d754cc0",
  1106 => x"87e0c302",
  1107 => x"1ed4f7c0",
  1108 => x"c70266c8",
  1109 => x"48a6cc87",
  1110 => x"87c578c0",
  1111 => x"c148a6cc",
  1112 => x"4966cc78",
  1113 => x"c487e2e5",
  1114 => x"487e7086",
  1115 => x"e8c20298",
  1116 => x"81cb4987",
  1117 => x"d0496997",
  1118 => x"d6c10299",
  1119 => x"fbc2c187",
  1120 => x"cb49744a",
  1121 => x"e6e4c191",
  1122 => x"c8797281",
  1123 => x"51ffc381",
  1124 => x"91de4974",
  1125 => x"4dc0ebc2",
  1126 => x"c1c28571",
  1127 => x"a5c17d97",
  1128 => x"51e0c049",
  1129 => x"97f2e5c2",
  1130 => x"87d202bf",
  1131 => x"a5c284c1",
  1132 => x"f2e5c24b",
  1133 => x"fe49db4a",
  1134 => x"c187ecfb",
  1135 => x"a5cd87db",
  1136 => x"c151c049",
  1137 => x"4ba5c284",
  1138 => x"49cb4a6e",
  1139 => x"87d7fbfe",
  1140 => x"c187c6c1",
  1141 => x"744af7c0",
  1142 => x"c191cb49",
  1143 => x"7281e6e4",
  1144 => x"f2e5c279",
  1145 => x"d802bf97",
  1146 => x"de497487",
  1147 => x"c284c191",
  1148 => x"714bc0eb",
  1149 => x"f2e5c283",
  1150 => x"fe49dd4a",
  1151 => x"d887e8fa",
  1152 => x"de4b7487",
  1153 => x"c0ebc293",
  1154 => x"49a3cb83",
  1155 => x"84c151c0",
  1156 => x"cb4a6e73",
  1157 => x"cefafe49",
  1158 => x"4866c487",
  1159 => x"a6c880c1",
  1160 => x"03acc758",
  1161 => x"6e87c5c0",
  1162 => x"87e0fc05",
  1163 => x"8ef44874",
  1164 => x"1e87fdf5",
  1165 => x"4b711e73",
  1166 => x"c191cb49",
  1167 => x"c881e6e4",
  1168 => x"e4c14aa1",
  1169 => x"501248d2",
  1170 => x"c04aa1c9",
  1171 => x"1248c1fa",
  1172 => x"c181ca50",
  1173 => x"1148d3e4",
  1174 => x"d3e4c150",
  1175 => x"1e49bf97",
  1176 => x"d2f649c0",
  1177 => x"d4eac287",
  1178 => x"c178de48",
  1179 => x"87dad749",
  1180 => x"87c0f526",
  1181 => x"494a711e",
  1182 => x"e4c191cb",
  1183 => x"81c881e6",
  1184 => x"eac24811",
  1185 => x"eac258d8",
  1186 => x"78c048ec",
  1187 => x"f9d649c1",
  1188 => x"1e4f2687",
  1189 => x"fac049c0",
  1190 => x"4f2687da",
  1191 => x"0299711e",
  1192 => x"e5c187d2",
  1193 => x"50c048fb",
  1194 => x"c9c180f7",
  1195 => x"e4c140f4",
  1196 => x"87ce78df",
  1197 => x"48f7e5c1",
  1198 => x"78d8e4c1",
  1199 => x"cac180fc",
  1200 => x"4f2678d3",
  1201 => x"5c5b5e0e",
  1202 => x"86f40e5d",
  1203 => x"cb494d71",
  1204 => x"e6e4c191",
  1205 => x"4aa1c881",
  1206 => x"c47ea1ca",
  1207 => x"eec248a6",
  1208 => x"6e78bfdc",
  1209 => x"c44bbf97",
  1210 => x"28734866",
  1211 => x"124c4b70",
  1212 => x"58a6cc48",
  1213 => x"84c19c70",
  1214 => x"699781c9",
  1215 => x"04acb749",
  1216 => x"4cc087c2",
  1217 => x"4abf976e",
  1218 => x"724966c8",
  1219 => x"c4b9ff31",
  1220 => x"48749966",
  1221 => x"4a703072",
  1222 => x"c2b07148",
  1223 => x"c058e0ee",
  1224 => x"c087ece4",
  1225 => x"87e2d449",
  1226 => x"f6c04975",
  1227 => x"8ef487e1",
  1228 => x"1e87fdf1",
  1229 => x"4b711e73",
  1230 => x"87c8fe49",
  1231 => x"c3fe4973",
  1232 => x"87f0f187",
  1233 => x"711e731e",
  1234 => x"4aa3c64b",
  1235 => x"c187db02",
  1236 => x"87d6028a",
  1237 => x"dac1028a",
  1238 => x"c0028a87",
  1239 => x"028a87fc",
  1240 => x"8a87e1c0",
  1241 => x"c187cb02",
  1242 => x"49c787db",
  1243 => x"c187c5fc",
  1244 => x"eac287de",
  1245 => x"c102bfec",
  1246 => x"c14887cb",
  1247 => x"f0eac288",
  1248 => x"87c1c158",
  1249 => x"bff0eac2",
  1250 => x"87f9c002",
  1251 => x"bfeceac2",
  1252 => x"c280c148",
  1253 => x"c058f0ea",
  1254 => x"eac287eb",
  1255 => x"c649bfec",
  1256 => x"f0eac289",
  1257 => x"a9b7c059",
  1258 => x"c287da03",
  1259 => x"c048ecea",
  1260 => x"c287d278",
  1261 => x"02bff0ea",
  1262 => x"eac287cb",
  1263 => x"c648bfec",
  1264 => x"f0eac280",
  1265 => x"d249c058",
  1266 => x"497387c0",
  1267 => x"87fff3c0",
  1268 => x"0e87e1ef",
  1269 => x"5d5c5b5e",
  1270 => x"86d0ff0e",
  1271 => x"c859a6dc",
  1272 => x"78c048a6",
  1273 => x"c4c180c4",
  1274 => x"80c47866",
  1275 => x"80c478c1",
  1276 => x"eac278c1",
  1277 => x"78c148f0",
  1278 => x"bfd4eac2",
  1279 => x"05a8de48",
  1280 => x"e0f387cb",
  1281 => x"cc497087",
  1282 => x"fccf59a6",
  1283 => x"87fde287",
  1284 => x"e287dfe3",
  1285 => x"4c7087ec",
  1286 => x"02acfbc0",
  1287 => x"d887fbc1",
  1288 => x"edc10566",
  1289 => x"66c0c187",
  1290 => x"6a82c44a",
  1291 => x"c11e727e",
  1292 => x"c448fee0",
  1293 => x"a1c84966",
  1294 => x"7141204a",
  1295 => x"87f905aa",
  1296 => x"4a265110",
  1297 => x"4866c0c1",
  1298 => x"78f3c8c1",
  1299 => x"81c7496a",
  1300 => x"c0c15174",
  1301 => x"81c84966",
  1302 => x"c0c151c1",
  1303 => x"81c94966",
  1304 => x"c0c151c0",
  1305 => x"81ca4966",
  1306 => x"1ec151c0",
  1307 => x"496a1ed8",
  1308 => x"d1e281c8",
  1309 => x"c186c887",
  1310 => x"c04866c4",
  1311 => x"87c701a8",
  1312 => x"c148a6c8",
  1313 => x"c187ce78",
  1314 => x"c14866c4",
  1315 => x"58a6d088",
  1316 => x"dde187c3",
  1317 => x"48a6d087",
  1318 => x"9c7478c2",
  1319 => x"87e5cd02",
  1320 => x"c14866c8",
  1321 => x"03a866c8",
  1322 => x"dc87dacd",
  1323 => x"78c048a6",
  1324 => x"78c080e8",
  1325 => x"7087cbe0",
  1326 => x"acd0c14c",
  1327 => x"87dac205",
  1328 => x"e27e66c4",
  1329 => x"497087ef",
  1330 => x"ff59a6c8",
  1331 => x"7087f3df",
  1332 => x"acecc04c",
  1333 => x"87edc105",
  1334 => x"cb4966c8",
  1335 => x"66c0c191",
  1336 => x"4aa1c481",
  1337 => x"a1c84d6a",
  1338 => x"5266c44a",
  1339 => x"79f4c9c1",
  1340 => x"87cedfff",
  1341 => x"029c4c70",
  1342 => x"fbc087d9",
  1343 => x"87d302ac",
  1344 => x"deff5574",
  1345 => x"4c7087fc",
  1346 => x"87c7029c",
  1347 => x"05acfbc0",
  1348 => x"c087edff",
  1349 => x"c1c255e0",
  1350 => x"7d97c055",
  1351 => x"6e4966d8",
  1352 => x"87db05a9",
  1353 => x"cc4866c8",
  1354 => x"ca04a866",
  1355 => x"4866c887",
  1356 => x"a6cc80c1",
  1357 => x"cc87c858",
  1358 => x"88c14866",
  1359 => x"ff58a6d0",
  1360 => x"7087ffdd",
  1361 => x"acd0c14c",
  1362 => x"d487c805",
  1363 => x"80c14866",
  1364 => x"c158a6d8",
  1365 => x"fd02acd0",
  1366 => x"e0c087e6",
  1367 => x"66d848a6",
  1368 => x"4866c478",
  1369 => x"a866e0c0",
  1370 => x"87ebc905",
  1371 => x"48a6e4c0",
  1372 => x"487478c0",
  1373 => x"7088fbc0",
  1374 => x"0298487e",
  1375 => x"4887edc9",
  1376 => x"7e7088cb",
  1377 => x"c1029848",
  1378 => x"c94887cd",
  1379 => x"487e7088",
  1380 => x"c1c40298",
  1381 => x"88c44887",
  1382 => x"98487e70",
  1383 => x"4887ce02",
  1384 => x"7e7088c1",
  1385 => x"c3029848",
  1386 => x"e1c887ec",
  1387 => x"48a6dc87",
  1388 => x"ff78f0c0",
  1389 => x"7087cbdc",
  1390 => x"acecc04c",
  1391 => x"87c4c002",
  1392 => x"5ca6e0c0",
  1393 => x"02acecc0",
  1394 => x"dbff87cd",
  1395 => x"4c7087f4",
  1396 => x"05acecc0",
  1397 => x"c087f3ff",
  1398 => x"c002acec",
  1399 => x"dbff87c4",
  1400 => x"1ec087e0",
  1401 => x"66d01eca",
  1402 => x"c191cb49",
  1403 => x"714866c8",
  1404 => x"58a6cc80",
  1405 => x"c44866c8",
  1406 => x"58a6d080",
  1407 => x"49bf66cc",
  1408 => x"87c2dcff",
  1409 => x"1ede1ec1",
  1410 => x"49bf66d4",
  1411 => x"87f6dbff",
  1412 => x"497086d0",
  1413 => x"c08909c0",
  1414 => x"c059a6ec",
  1415 => x"c04866e8",
  1416 => x"eec006a8",
  1417 => x"66e8c087",
  1418 => x"03a8dd48",
  1419 => x"c487e4c0",
  1420 => x"c049bf66",
  1421 => x"c08166e8",
  1422 => x"e8c051e0",
  1423 => x"81c14966",
  1424 => x"81bf66c4",
  1425 => x"c051c1c2",
  1426 => x"c24966e8",
  1427 => x"bf66c481",
  1428 => x"6e51c081",
  1429 => x"f3c8c148",
  1430 => x"c8496e78",
  1431 => x"5166d081",
  1432 => x"81c9496e",
  1433 => x"6e5166d4",
  1434 => x"dc81ca49",
  1435 => x"66d05166",
  1436 => x"d480c148",
  1437 => x"66c858a6",
  1438 => x"a866cc48",
  1439 => x"87cbc004",
  1440 => x"c14866c8",
  1441 => x"58a6cc80",
  1442 => x"cc87e1c5",
  1443 => x"88c14866",
  1444 => x"c558a6d0",
  1445 => x"dbff87d6",
  1446 => x"497087db",
  1447 => x"59a6ecc0",
  1448 => x"87d1dbff",
  1449 => x"e0c04970",
  1450 => x"66dc59a6",
  1451 => x"a8ecc048",
  1452 => x"87cac005",
  1453 => x"c048a6dc",
  1454 => x"c07866e8",
  1455 => x"d8ff87c4",
  1456 => x"66c887c0",
  1457 => x"c191cb49",
  1458 => x"714866c0",
  1459 => x"4a7e7080",
  1460 => x"496e82c8",
  1461 => x"e8c081ca",
  1462 => x"66dc5166",
  1463 => x"c081c149",
  1464 => x"c18966e8",
  1465 => x"70307148",
  1466 => x"7189c149",
  1467 => x"eec27a97",
  1468 => x"c049bfdc",
  1469 => x"972966e8",
  1470 => x"71484a6a",
  1471 => x"a6f0c098",
  1472 => x"c4496e58",
  1473 => x"c04d6981",
  1474 => x"c44866e0",
  1475 => x"c002a866",
  1476 => x"a6c487c8",
  1477 => x"c078c048",
  1478 => x"a6c487c5",
  1479 => x"c478c148",
  1480 => x"e0c01e66",
  1481 => x"ff49751e",
  1482 => x"c887dbd7",
  1483 => x"c04c7086",
  1484 => x"c106acb7",
  1485 => x"857487d4",
  1486 => x"7449e0c0",
  1487 => x"c14b7589",
  1488 => x"714ac7e1",
  1489 => x"87dfe5fe",
  1490 => x"e4c085c2",
  1491 => x"80c14866",
  1492 => x"58a6e8c0",
  1493 => x"4966ecc0",
  1494 => x"a97081c1",
  1495 => x"87c8c002",
  1496 => x"c048a6c4",
  1497 => x"87c5c078",
  1498 => x"c148a6c4",
  1499 => x"1e66c478",
  1500 => x"c049a4c2",
  1501 => x"887148e0",
  1502 => x"751e4970",
  1503 => x"c5d6ff49",
  1504 => x"c086c887",
  1505 => x"ff01a8b7",
  1506 => x"e4c087c0",
  1507 => x"d1c00266",
  1508 => x"c9496e87",
  1509 => x"66e4c081",
  1510 => x"c1486e51",
  1511 => x"c078c4cb",
  1512 => x"496e87cc",
  1513 => x"51c281c9",
  1514 => x"ccc1486e",
  1515 => x"66c878f3",
  1516 => x"a866cc48",
  1517 => x"87cbc004",
  1518 => x"c14866c8",
  1519 => x"58a6cc80",
  1520 => x"cc87e9c0",
  1521 => x"88c14866",
  1522 => x"c058a6d0",
  1523 => x"d4ff87de",
  1524 => x"4c7087e0",
  1525 => x"c187d5c0",
  1526 => x"c005acc6",
  1527 => x"66d087c8",
  1528 => x"d480c148",
  1529 => x"d4ff58a6",
  1530 => x"4c7087c8",
  1531 => x"c14866d4",
  1532 => x"58a6d880",
  1533 => x"c0029c74",
  1534 => x"66c887cb",
  1535 => x"66c8c148",
  1536 => x"e6f204a8",
  1537 => x"e0d3ff87",
  1538 => x"4866c887",
  1539 => x"c003a8c7",
  1540 => x"eac287e5",
  1541 => x"78c048f0",
  1542 => x"cb4966c8",
  1543 => x"66c0c191",
  1544 => x"4aa1c481",
  1545 => x"52c04a6a",
  1546 => x"4866c879",
  1547 => x"a6cc80c1",
  1548 => x"04a8c758",
  1549 => x"ff87dbff",
  1550 => x"ddff8ed0",
  1551 => x"6f4c87f2",
  1552 => x"2a206461",
  1553 => x"3a00202e",
  1554 => x"731e0020",
  1555 => x"9b4b711e",
  1556 => x"c287c602",
  1557 => x"c048ecea",
  1558 => x"c21ec778",
  1559 => x"49bfecea",
  1560 => x"e6e4c11e",
  1561 => x"d4eac21e",
  1562 => x"e6ed49bf",
  1563 => x"c286cc87",
  1564 => x"49bfd4ea",
  1565 => x"7387e5e8",
  1566 => x"87c8029b",
  1567 => x"49e6e4c1",
  1568 => x"87dde2c0",
  1569 => x"87ecdcff",
  1570 => x"87d4c71e",
  1571 => x"f9fe49c1",
  1572 => x"fae8fe87",
  1573 => x"02987087",
  1574 => x"f1fe87cd",
  1575 => x"987087f5",
  1576 => x"c187c402",
  1577 => x"c087c24a",
  1578 => x"059a724a",
  1579 => x"1ec087ce",
  1580 => x"49d9e3c1",
  1581 => x"87d6efc0",
  1582 => x"87fe86c4",
  1583 => x"e3c11ec0",
  1584 => x"efc049e4",
  1585 => x"1ec087c8",
  1586 => x"87def8c0",
  1587 => x"eec04970",
  1588 => x"cac387fc",
  1589 => x"268ef887",
  1590 => x"2044534f",
  1591 => x"6c696166",
  1592 => x"002e6465",
  1593 => x"746f6f42",
  1594 => x"2e676e69",
  1595 => x"1e002e2e",
  1596 => x"87ebe5c0",
  1597 => x"87e1f2c0",
  1598 => x"4f2687f6",
  1599 => x"eceac21e",
  1600 => x"c278c048",
  1601 => x"c048d4ea",
  1602 => x"87fcfd78",
  1603 => x"48c087e1",
  1604 => x"00004f26",
  1605 => x"00000001",
  1606 => x"78452080",
  1607 => x"80007469",
  1608 => x"63614220",
  1609 => x"1037006b",
  1610 => x"2ac00000",
  1611 => x"00000000",
  1612 => x"00103700",
  1613 => x"002ade00",
  1614 => x"00000000",
  1615 => x"00001037",
  1616 => x"00002afc",
  1617 => x"37000000",
  1618 => x"1a000010",
  1619 => x"0000002b",
  1620 => x"10370000",
  1621 => x"2b380000",
  1622 => x"00000000",
  1623 => x"00103700",
  1624 => x"002b5600",
  1625 => x"00000000",
  1626 => x"00001037",
  1627 => x"00002b74",
  1628 => x"74000000",
  1629 => x"00000012",
  1630 => x"00000000",
  1631 => x"13440000",
  1632 => x"00000000",
  1633 => x"00000000",
  1634 => x"f0fe1e00",
  1635 => x"cd78c048",
  1636 => x"26097909",
  1637 => x"fe1e1e4f",
  1638 => x"487ebff0",
  1639 => x"1e4f2626",
  1640 => x"c148f0fe",
  1641 => x"1e4f2678",
  1642 => x"c048f0fe",
  1643 => x"1e4f2678",
  1644 => x"52c04a71",
  1645 => x"0e4f2652",
  1646 => x"5d5c5b5e",
  1647 => x"7186f40e",
  1648 => x"7e6d974d",
  1649 => x"974ca5c1",
  1650 => x"a6c8486c",
  1651 => x"c4486e58",
  1652 => x"c505a866",
  1653 => x"c048ff87",
  1654 => x"caff87e6",
  1655 => x"49a5c287",
  1656 => x"714b6c97",
  1657 => x"6b974ba3",
  1658 => x"7e6c974b",
  1659 => x"80c1486e",
  1660 => x"c758a6c8",
  1661 => x"58a6cc98",
  1662 => x"fe7c9770",
  1663 => x"487387e1",
  1664 => x"4d268ef4",
  1665 => x"4b264c26",
  1666 => x"5e0e4f26",
  1667 => x"f40e5c5b",
  1668 => x"d84c7186",
  1669 => x"ffc34a66",
  1670 => x"4ba4c29a",
  1671 => x"73496c97",
  1672 => x"517249a1",
  1673 => x"6e7e6c97",
  1674 => x"c880c148",
  1675 => x"98c758a6",
  1676 => x"7058a6cc",
  1677 => x"ff8ef454",
  1678 => x"1e1e87ca",
  1679 => x"e087e8fd",
  1680 => x"c0494abf",
  1681 => x"0299c0e0",
  1682 => x"1e7287cb",
  1683 => x"49d2eec2",
  1684 => x"c487f7fe",
  1685 => x"87fdfc86",
  1686 => x"c2fd7e70",
  1687 => x"4f262687",
  1688 => x"d2eec21e",
  1689 => x"87c7fd49",
  1690 => x"49fae8c1",
  1691 => x"c387dafc",
  1692 => x"4f2687f7",
  1693 => x"5c5b5e0e",
  1694 => x"4d710e5d",
  1695 => x"49d2eec2",
  1696 => x"7087f4fc",
  1697 => x"abb7c04b",
  1698 => x"87c2c304",
  1699 => x"05abf0c3",
  1700 => x"edc187c9",
  1701 => x"78c148d8",
  1702 => x"c387e3c2",
  1703 => x"c905abe0",
  1704 => x"dcedc187",
  1705 => x"c278c148",
  1706 => x"edc187d4",
  1707 => x"c602bfdc",
  1708 => x"a3c0c287",
  1709 => x"7387c24c",
  1710 => x"d8edc14c",
  1711 => x"e0c002bf",
  1712 => x"c4497487",
  1713 => x"c19129b7",
  1714 => x"7481f8ee",
  1715 => x"c29acf4a",
  1716 => x"7248c192",
  1717 => x"ff4a7030",
  1718 => x"694872ba",
  1719 => x"db797098",
  1720 => x"c4497487",
  1721 => x"c19129b7",
  1722 => x"7481f8ee",
  1723 => x"c29acf4a",
  1724 => x"7248c392",
  1725 => x"484a7030",
  1726 => x"7970b069",
  1727 => x"c0059d75",
  1728 => x"d0ff87f0",
  1729 => x"78e1c848",
  1730 => x"c548d4ff",
  1731 => x"dcedc178",
  1732 => x"87c302bf",
  1733 => x"c178e0c3",
  1734 => x"02bfd8ed",
  1735 => x"d4ff87c6",
  1736 => x"78f0c348",
  1737 => x"7348d4ff",
  1738 => x"48d0ff78",
  1739 => x"c078e1c8",
  1740 => x"edc178e0",
  1741 => x"78c048dc",
  1742 => x"48d8edc1",
  1743 => x"eec278c0",
  1744 => x"f2f949d2",
  1745 => x"c04b7087",
  1746 => x"fc03abb7",
  1747 => x"48c087fe",
  1748 => x"4c264d26",
  1749 => x"4f264b26",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"494a711e",
  1753 => x"2687cdfc",
  1754 => x"4ac01e4f",
  1755 => x"91c44972",
  1756 => x"81f8eec1",
  1757 => x"82c179c0",
  1758 => x"04aab7d0",
  1759 => x"4f2687ee",
  1760 => x"5c5b5e0e",
  1761 => x"4d710e5d",
  1762 => x"7587dcf8",
  1763 => x"2ab7c44a",
  1764 => x"f8eec192",
  1765 => x"cf4c7582",
  1766 => x"6a94c29c",
  1767 => x"2b744b49",
  1768 => x"48c29bc3",
  1769 => x"4c703074",
  1770 => x"4874bcff",
  1771 => x"7a709871",
  1772 => x"7387ecf7",
  1773 => x"87d8fe48",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"48d0ff1e",
  1791 => x"7178e1c8",
  1792 => x"08d4ff48",
  1793 => x"1e4f2678",
  1794 => x"c848d0ff",
  1795 => x"487178e1",
  1796 => x"7808d4ff",
  1797 => x"ff4866c4",
  1798 => x"267808d4",
  1799 => x"4a711e4f",
  1800 => x"1e4966c4",
  1801 => x"deff4972",
  1802 => x"48d0ff87",
  1803 => x"2678e0c0",
  1804 => x"731e4f26",
  1805 => x"c84b711e",
  1806 => x"731e4966",
  1807 => x"a2e0c14a",
  1808 => x"87d9ff49",
  1809 => x"2687c426",
  1810 => x"264c264d",
  1811 => x"1e4f264b",
  1812 => x"c34ad4ff",
  1813 => x"d0ff7aff",
  1814 => x"78e1c048",
  1815 => x"eec27ade",
  1816 => x"497abfdc",
  1817 => x"7028c848",
  1818 => x"d048717a",
  1819 => x"717a7028",
  1820 => x"7028d848",
  1821 => x"48d0ff7a",
  1822 => x"2678e0c0",
  1823 => x"d0ff1e4f",
  1824 => x"78c9c848",
  1825 => x"d4ff4871",
  1826 => x"4f267808",
  1827 => x"494a711e",
  1828 => x"d0ff87eb",
  1829 => x"2678c848",
  1830 => x"1e731e4f",
  1831 => x"eec24b71",
  1832 => x"c302bfec",
  1833 => x"87ebc287",
  1834 => x"c848d0ff",
  1835 => x"497378c9",
  1836 => x"ffb1e0c0",
  1837 => x"787148d4",
  1838 => x"48e0eec2",
  1839 => x"66c878c0",
  1840 => x"c387c502",
  1841 => x"87c249ff",
  1842 => x"eec249c0",
  1843 => x"66cc59e8",
  1844 => x"c587c602",
  1845 => x"c44ad5d5",
  1846 => x"ffffcf87",
  1847 => x"eceec24a",
  1848 => x"eceec25a",
  1849 => x"c478c148",
  1850 => x"264d2687",
  1851 => x"264b264c",
  1852 => x"5b5e0e4f",
  1853 => x"710e5d5c",
  1854 => x"e8eec24a",
  1855 => x"9a724cbf",
  1856 => x"4987cb02",
  1857 => x"f2c191c8",
  1858 => x"83714bcf",
  1859 => x"f6c187c4",
  1860 => x"4dc04bcf",
  1861 => x"99744913",
  1862 => x"bfe4eec2",
  1863 => x"48d4ffb9",
  1864 => x"b7c17871",
  1865 => x"b7c8852c",
  1866 => x"87e804ad",
  1867 => x"bfe0eec2",
  1868 => x"c280c848",
  1869 => x"fe58e4ee",
  1870 => x"731e87ef",
  1871 => x"134b711e",
  1872 => x"cb029a4a",
  1873 => x"fe497287",
  1874 => x"4a1387e7",
  1875 => x"87f5059a",
  1876 => x"1e87dafe",
  1877 => x"bfe0eec2",
  1878 => x"e0eec249",
  1879 => x"78a1c148",
  1880 => x"a9b7c0c4",
  1881 => x"ff87db03",
  1882 => x"eec248d4",
  1883 => x"c278bfe4",
  1884 => x"49bfe0ee",
  1885 => x"48e0eec2",
  1886 => x"c478a1c1",
  1887 => x"04a9b7c0",
  1888 => x"d0ff87e5",
  1889 => x"c278c848",
  1890 => x"c048ecee",
  1891 => x"004f2678",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"5f5f0000",
  1895 => x"00000000",
  1896 => x"03000303",
  1897 => x"14000003",
  1898 => x"7f147f7f",
  1899 => x"0000147f",
  1900 => x"6b6b2e24",
  1901 => x"4c00123a",
  1902 => x"6c18366a",
  1903 => x"30003256",
  1904 => x"77594f7e",
  1905 => x"0040683a",
  1906 => x"03070400",
  1907 => x"00000000",
  1908 => x"633e1c00",
  1909 => x"00000041",
  1910 => x"3e634100",
  1911 => x"0800001c",
  1912 => x"1c1c3e2a",
  1913 => x"00082a3e",
  1914 => x"3e3e0808",
  1915 => x"00000808",
  1916 => x"60e08000",
  1917 => x"00000000",
  1918 => x"08080808",
  1919 => x"00000808",
  1920 => x"60600000",
  1921 => x"40000000",
  1922 => x"0c183060",
  1923 => x"00010306",
  1924 => x"4d597f3e",
  1925 => x"00003e7f",
  1926 => x"7f7f0604",
  1927 => x"00000000",
  1928 => x"59716342",
  1929 => x"0000464f",
  1930 => x"49496322",
  1931 => x"1800367f",
  1932 => x"7f13161c",
  1933 => x"0000107f",
  1934 => x"45456727",
  1935 => x"0000397d",
  1936 => x"494b7e3c",
  1937 => x"00003079",
  1938 => x"79710101",
  1939 => x"0000070f",
  1940 => x"49497f36",
  1941 => x"0000367f",
  1942 => x"69494f06",
  1943 => x"00001e3f",
  1944 => x"66660000",
  1945 => x"00000000",
  1946 => x"66e68000",
  1947 => x"00000000",
  1948 => x"14140808",
  1949 => x"00002222",
  1950 => x"14141414",
  1951 => x"00001414",
  1952 => x"14142222",
  1953 => x"00000808",
  1954 => x"59510302",
  1955 => x"3e00060f",
  1956 => x"555d417f",
  1957 => x"00001e1f",
  1958 => x"09097f7e",
  1959 => x"00007e7f",
  1960 => x"49497f7f",
  1961 => x"0000367f",
  1962 => x"41633e1c",
  1963 => x"00004141",
  1964 => x"63417f7f",
  1965 => x"00001c3e",
  1966 => x"49497f7f",
  1967 => x"00004141",
  1968 => x"09097f7f",
  1969 => x"00000101",
  1970 => x"49417f3e",
  1971 => x"00007a7b",
  1972 => x"08087f7f",
  1973 => x"00007f7f",
  1974 => x"7f7f4100",
  1975 => x"00000041",
  1976 => x"40406020",
  1977 => x"7f003f7f",
  1978 => x"361c087f",
  1979 => x"00004163",
  1980 => x"40407f7f",
  1981 => x"7f004040",
  1982 => x"060c067f",
  1983 => x"7f007f7f",
  1984 => x"180c067f",
  1985 => x"00007f7f",
  1986 => x"41417f3e",
  1987 => x"00003e7f",
  1988 => x"09097f7f",
  1989 => x"3e00060f",
  1990 => x"7f61417f",
  1991 => x"0000407e",
  1992 => x"19097f7f",
  1993 => x"0000667f",
  1994 => x"594d6f26",
  1995 => x"0000327b",
  1996 => x"7f7f0101",
  1997 => x"00000101",
  1998 => x"40407f3f",
  1999 => x"00003f7f",
  2000 => x"70703f0f",
  2001 => x"7f000f3f",
  2002 => x"3018307f",
  2003 => x"41007f7f",
  2004 => x"1c1c3663",
  2005 => x"01416336",
  2006 => x"7c7c0603",
  2007 => x"61010306",
  2008 => x"474d5971",
  2009 => x"00004143",
  2010 => x"417f7f00",
  2011 => x"01000041",
  2012 => x"180c0603",
  2013 => x"00406030",
  2014 => x"7f414100",
  2015 => x"0800007f",
  2016 => x"0603060c",
  2017 => x"8000080c",
  2018 => x"80808080",
  2019 => x"00008080",
  2020 => x"07030000",
  2021 => x"00000004",
  2022 => x"54547420",
  2023 => x"0000787c",
  2024 => x"44447f7f",
  2025 => x"0000387c",
  2026 => x"44447c38",
  2027 => x"00000044",
  2028 => x"44447c38",
  2029 => x"00007f7f",
  2030 => x"54547c38",
  2031 => x"0000185c",
  2032 => x"057f7e04",
  2033 => x"00000005",
  2034 => x"a4a4bc18",
  2035 => x"00007cfc",
  2036 => x"04047f7f",
  2037 => x"0000787c",
  2038 => x"7d3d0000",
  2039 => x"00000040",
  2040 => x"fd808080",
  2041 => x"0000007d",
  2042 => x"38107f7f",
  2043 => x"0000446c",
  2044 => x"7f3f0000",
  2045 => x"7c000040",
  2046 => x"0c180c7c",
  2047 => x"0000787c",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
