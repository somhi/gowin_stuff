
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"04",x"7c",x"7c"),
     1 => (x"00",x"00",x"78",x"7c"),
     2 => (x"44",x"44",x"7c",x"38"),
     3 => (x"00",x"00",x"38",x"7c"),
     4 => (x"24",x"24",x"fc",x"fc"),
     5 => (x"00",x"00",x"18",x"3c"),
     6 => (x"24",x"24",x"3c",x"18"),
     7 => (x"00",x"00",x"fc",x"fc"),
     8 => (x"04",x"04",x"7c",x"7c"),
     9 => (x"00",x"00",x"08",x"0c"),
    10 => (x"54",x"54",x"5c",x"48"),
    11 => (x"00",x"00",x"20",x"74"),
    12 => (x"44",x"7f",x"3f",x"04"),
    13 => (x"00",x"00",x"00",x"44"),
    14 => (x"40",x"40",x"7c",x"3c"),
    15 => (x"00",x"00",x"7c",x"7c"),
    16 => (x"60",x"60",x"3c",x"1c"),
    17 => (x"3c",x"00",x"1c",x"3c"),
    18 => (x"60",x"30",x"60",x"7c"),
    19 => (x"44",x"00",x"3c",x"7c"),
    20 => (x"38",x"10",x"38",x"6c"),
    21 => (x"00",x"00",x"44",x"6c"),
    22 => (x"60",x"e0",x"bc",x"1c"),
    23 => (x"00",x"00",x"1c",x"3c"),
    24 => (x"5c",x"74",x"64",x"44"),
    25 => (x"00",x"00",x"44",x"4c"),
    26 => (x"77",x"3e",x"08",x"08"),
    27 => (x"00",x"00",x"41",x"41"),
    28 => (x"7f",x"7f",x"00",x"00"),
    29 => (x"00",x"00",x"00",x"00"),
    30 => (x"3e",x"77",x"41",x"41"),
    31 => (x"02",x"00",x"08",x"08"),
    32 => (x"02",x"03",x"01",x"01"),
    33 => (x"7f",x"00",x"01",x"02"),
    34 => (x"7f",x"7f",x"7f",x"7f"),
    35 => (x"08",x"00",x"7f",x"7f"),
    36 => (x"3e",x"1c",x"1c",x"08"),
    37 => (x"7f",x"7f",x"7f",x"3e"),
    38 => (x"1c",x"3e",x"3e",x"7f"),
    39 => (x"00",x"08",x"08",x"1c"),
    40 => (x"7c",x"7c",x"18",x"10"),
    41 => (x"00",x"00",x"10",x"18"),
    42 => (x"7c",x"7c",x"30",x"10"),
    43 => (x"10",x"00",x"10",x"30"),
    44 => (x"78",x"60",x"60",x"30"),
    45 => (x"42",x"00",x"06",x"1e"),
    46 => (x"3c",x"18",x"3c",x"66"),
    47 => (x"78",x"00",x"42",x"66"),
    48 => (x"c6",x"c2",x"6a",x"38"),
    49 => (x"60",x"00",x"38",x"6c"),
    50 => (x"00",x"60",x"00",x"00"),
    51 => (x"0e",x"00",x"60",x"00"),
    52 => (x"5d",x"5c",x"5b",x"5e"),
    53 => (x"4c",x"71",x"1e",x"0e"),
    54 => (x"bf",x"fd",x"ee",x"c2"),
    55 => (x"c0",x"4b",x"c0",x"4d"),
    56 => (x"02",x"ab",x"74",x"1e"),
    57 => (x"a6",x"c4",x"87",x"c7"),
    58 => (x"c5",x"78",x"c0",x"48"),
    59 => (x"48",x"a6",x"c4",x"87"),
    60 => (x"66",x"c4",x"78",x"c1"),
    61 => (x"ee",x"49",x"73",x"1e"),
    62 => (x"86",x"c8",x"87",x"df"),
    63 => (x"ef",x"49",x"e0",x"c0"),
    64 => (x"a5",x"c4",x"87",x"ef"),
    65 => (x"f0",x"49",x"6a",x"4a"),
    66 => (x"c6",x"f1",x"87",x"f0"),
    67 => (x"c1",x"85",x"cb",x"87"),
    68 => (x"ab",x"b7",x"c8",x"83"),
    69 => (x"87",x"c7",x"ff",x"04"),
    70 => (x"26",x"4d",x"26",x"26"),
    71 => (x"26",x"4b",x"26",x"4c"),
    72 => (x"4a",x"71",x"1e",x"4f"),
    73 => (x"5a",x"c1",x"ef",x"c2"),
    74 => (x"48",x"c1",x"ef",x"c2"),
    75 => (x"fe",x"49",x"78",x"c7"),
    76 => (x"4f",x"26",x"87",x"dd"),
    77 => (x"71",x"1e",x"73",x"1e"),
    78 => (x"aa",x"b7",x"c0",x"4a"),
    79 => (x"c2",x"87",x"d3",x"03"),
    80 => (x"05",x"bf",x"f8",x"d3"),
    81 => (x"4b",x"c1",x"87",x"c4"),
    82 => (x"4b",x"c0",x"87",x"c2"),
    83 => (x"5b",x"fc",x"d3",x"c2"),
    84 => (x"d3",x"c2",x"87",x"c4"),
    85 => (x"d3",x"c2",x"5a",x"fc"),
    86 => (x"c1",x"4a",x"bf",x"f8"),
    87 => (x"a2",x"c0",x"c1",x"9a"),
    88 => (x"87",x"e8",x"ec",x"49"),
    89 => (x"d3",x"c2",x"48",x"fc"),
    90 => (x"fe",x"78",x"bf",x"f8"),
    91 => (x"71",x"1e",x"87",x"ef"),
    92 => (x"1e",x"66",x"c4",x"4a"),
    93 => (x"f9",x"ea",x"49",x"72"),
    94 => (x"4f",x"26",x"26",x"87"),
    95 => (x"ff",x"4a",x"71",x"1e"),
    96 => (x"ff",x"c3",x"48",x"d4"),
    97 => (x"48",x"d0",x"ff",x"78"),
    98 => (x"ff",x"78",x"e1",x"c0"),
    99 => (x"78",x"c1",x"48",x"d4"),
   100 => (x"31",x"c4",x"49",x"72"),
   101 => (x"d0",x"ff",x"78",x"71"),
   102 => (x"78",x"e0",x"c0",x"48"),
   103 => (x"c2",x"1e",x"4f",x"26"),
   104 => (x"49",x"bf",x"f8",x"d3"),
   105 => (x"c2",x"87",x"f9",x"e6"),
   106 => (x"e8",x"48",x"f5",x"ee"),
   107 => (x"ee",x"c2",x"78",x"bf"),
   108 => (x"bf",x"ec",x"48",x"f1"),
   109 => (x"f5",x"ee",x"c2",x"78"),
   110 => (x"c3",x"49",x"4a",x"bf"),
   111 => (x"b7",x"c8",x"99",x"ff"),
   112 => (x"71",x"48",x"72",x"2a"),
   113 => (x"fd",x"ee",x"c2",x"b0"),
   114 => (x"0e",x"4f",x"26",x"58"),
   115 => (x"5d",x"5c",x"5b",x"5e"),
   116 => (x"ff",x"4b",x"71",x"0e"),
   117 => (x"ee",x"c2",x"87",x"c8"),
   118 => (x"50",x"c0",x"48",x"f0"),
   119 => (x"df",x"e6",x"49",x"73"),
   120 => (x"4c",x"49",x"70",x"87"),
   121 => (x"ee",x"cb",x"9c",x"c2"),
   122 => (x"87",x"d4",x"cc",x"49"),
   123 => (x"c2",x"4d",x"49",x"70"),
   124 => (x"bf",x"97",x"f0",x"ee"),
   125 => (x"87",x"e2",x"c1",x"05"),
   126 => (x"c2",x"49",x"66",x"d0"),
   127 => (x"99",x"bf",x"f9",x"ee"),
   128 => (x"d4",x"87",x"d6",x"05"),
   129 => (x"ee",x"c2",x"49",x"66"),
   130 => (x"05",x"99",x"bf",x"f1"),
   131 => (x"49",x"73",x"87",x"cb"),
   132 => (x"70",x"87",x"ed",x"e5"),
   133 => (x"c1",x"c1",x"02",x"98"),
   134 => (x"fe",x"4c",x"c1",x"87"),
   135 => (x"49",x"75",x"87",x"c0"),
   136 => (x"70",x"87",x"e9",x"cb"),
   137 => (x"87",x"c6",x"02",x"98"),
   138 => (x"48",x"f0",x"ee",x"c2"),
   139 => (x"ee",x"c2",x"50",x"c1"),
   140 => (x"05",x"bf",x"97",x"f0"),
   141 => (x"c2",x"87",x"e3",x"c0"),
   142 => (x"49",x"bf",x"f9",x"ee"),
   143 => (x"05",x"99",x"66",x"d0"),
   144 => (x"c2",x"87",x"d6",x"ff"),
   145 => (x"49",x"bf",x"f1",x"ee"),
   146 => (x"05",x"99",x"66",x"d4"),
   147 => (x"73",x"87",x"ca",x"ff"),
   148 => (x"87",x"ec",x"e4",x"49"),
   149 => (x"fe",x"05",x"98",x"70"),
   150 => (x"48",x"74",x"87",x"ff"),
   151 => (x"0e",x"87",x"fa",x"fa"),
   152 => (x"5d",x"5c",x"5b",x"5e"),
   153 => (x"c0",x"86",x"f8",x"0e"),
   154 => (x"bf",x"ec",x"4c",x"4d"),
   155 => (x"48",x"a6",x"c4",x"7e"),
   156 => (x"bf",x"fd",x"ee",x"c2"),
   157 => (x"c0",x"1e",x"c1",x"78"),
   158 => (x"fd",x"49",x"c7",x"1e"),
   159 => (x"86",x"c8",x"87",x"cd"),
   160 => (x"cd",x"02",x"98",x"70"),
   161 => (x"fa",x"49",x"ff",x"87"),
   162 => (x"da",x"c1",x"87",x"ea"),
   163 => (x"87",x"f0",x"e3",x"49"),
   164 => (x"ee",x"c2",x"4d",x"c1"),
   165 => (x"02",x"bf",x"97",x"f0"),
   166 => (x"d3",x"c2",x"87",x"cf"),
   167 => (x"c1",x"49",x"bf",x"e0"),
   168 => (x"e4",x"d3",x"c2",x"b9"),
   169 => (x"d3",x"fb",x"71",x"59"),
   170 => (x"f5",x"ee",x"c2",x"87"),
   171 => (x"d3",x"c2",x"4b",x"bf"),
   172 => (x"c1",x"05",x"bf",x"f8"),
   173 => (x"a6",x"c4",x"87",x"d9"),
   174 => (x"c0",x"c0",x"c8",x"48"),
   175 => (x"e4",x"d3",x"c2",x"78"),
   176 => (x"bf",x"97",x"6e",x"7e"),
   177 => (x"c1",x"48",x"6e",x"49"),
   178 => (x"71",x"7e",x"70",x"80"),
   179 => (x"70",x"87",x"f1",x"e2"),
   180 => (x"87",x"c3",x"02",x"98"),
   181 => (x"c4",x"b3",x"66",x"c4"),
   182 => (x"b7",x"c1",x"48",x"66"),
   183 => (x"58",x"a6",x"c8",x"28"),
   184 => (x"ff",x"05",x"98",x"70"),
   185 => (x"fd",x"c3",x"87",x"db"),
   186 => (x"87",x"d4",x"e2",x"49"),
   187 => (x"e2",x"49",x"fa",x"c3"),
   188 => (x"49",x"73",x"87",x"ce"),
   189 => (x"71",x"99",x"ff",x"c3"),
   190 => (x"f9",x"49",x"c0",x"1e"),
   191 => (x"49",x"73",x"87",x"f0"),
   192 => (x"71",x"29",x"b7",x"c8"),
   193 => (x"f9",x"49",x"c1",x"1e"),
   194 => (x"86",x"c8",x"87",x"e4"),
   195 => (x"c2",x"87",x"fa",x"c5"),
   196 => (x"4b",x"bf",x"f9",x"ee"),
   197 => (x"87",x"dd",x"02",x"9b"),
   198 => (x"bf",x"f4",x"d3",x"c2"),
   199 => (x"87",x"ec",x"c7",x"49"),
   200 => (x"c4",x"05",x"98",x"70"),
   201 => (x"d2",x"4b",x"c0",x"87"),
   202 => (x"49",x"e0",x"c2",x"87"),
   203 => (x"c2",x"87",x"d1",x"c7"),
   204 => (x"c6",x"58",x"f8",x"d3"),
   205 => (x"f4",x"d3",x"c2",x"87"),
   206 => (x"73",x"78",x"c0",x"48"),
   207 => (x"05",x"99",x"c2",x"49"),
   208 => (x"eb",x"c3",x"87",x"ce"),
   209 => (x"87",x"f8",x"e0",x"49"),
   210 => (x"99",x"c2",x"49",x"70"),
   211 => (x"87",x"c2",x"c0",x"02"),
   212 => (x"49",x"73",x"4c",x"fb"),
   213 => (x"ce",x"05",x"99",x"c1"),
   214 => (x"49",x"f4",x"c3",x"87"),
   215 => (x"70",x"87",x"e1",x"e0"),
   216 => (x"02",x"99",x"c2",x"49"),
   217 => (x"fa",x"87",x"c2",x"c0"),
   218 => (x"c8",x"49",x"73",x"4c"),
   219 => (x"87",x"cd",x"05",x"99"),
   220 => (x"e0",x"49",x"f5",x"c3"),
   221 => (x"49",x"70",x"87",x"ca"),
   222 => (x"d6",x"02",x"99",x"c2"),
   223 => (x"c1",x"ef",x"c2",x"87"),
   224 => (x"ca",x"c0",x"02",x"bf"),
   225 => (x"88",x"c1",x"48",x"87"),
   226 => (x"58",x"c5",x"ef",x"c2"),
   227 => (x"ff",x"87",x"c2",x"c0"),
   228 => (x"73",x"4d",x"c1",x"4c"),
   229 => (x"05",x"99",x"c4",x"49"),
   230 => (x"c3",x"87",x"ce",x"c0"),
   231 => (x"df",x"ff",x"49",x"f2"),
   232 => (x"49",x"70",x"87",x"de"),
   233 => (x"dc",x"02",x"99",x"c2"),
   234 => (x"c1",x"ef",x"c2",x"87"),
   235 => (x"c7",x"48",x"7e",x"bf"),
   236 => (x"c0",x"03",x"a8",x"b7"),
   237 => (x"48",x"6e",x"87",x"cb"),
   238 => (x"ef",x"c2",x"80",x"c1"),
   239 => (x"c2",x"c0",x"58",x"c5"),
   240 => (x"c1",x"4c",x"fe",x"87"),
   241 => (x"49",x"fd",x"c3",x"4d"),
   242 => (x"87",x"f4",x"de",x"ff"),
   243 => (x"99",x"c2",x"49",x"70"),
   244 => (x"87",x"d5",x"c0",x"02"),
   245 => (x"bf",x"c1",x"ef",x"c2"),
   246 => (x"87",x"c9",x"c0",x"02"),
   247 => (x"48",x"c1",x"ef",x"c2"),
   248 => (x"c2",x"c0",x"78",x"c0"),
   249 => (x"c1",x"4c",x"fd",x"87"),
   250 => (x"49",x"fa",x"c3",x"4d"),
   251 => (x"87",x"d0",x"de",x"ff"),
   252 => (x"99",x"c2",x"49",x"70"),
   253 => (x"87",x"d9",x"c0",x"02"),
   254 => (x"bf",x"c1",x"ef",x"c2"),
   255 => (x"a8",x"b7",x"c7",x"48"),
   256 => (x"87",x"c9",x"c0",x"03"),
   257 => (x"48",x"c1",x"ef",x"c2"),
   258 => (x"c2",x"c0",x"78",x"c7"),
   259 => (x"c1",x"4c",x"fc",x"87"),
   260 => (x"ac",x"b7",x"c0",x"4d"),
   261 => (x"87",x"d3",x"c0",x"03"),
   262 => (x"c1",x"48",x"66",x"c4"),
   263 => (x"7e",x"70",x"80",x"d8"),
   264 => (x"c0",x"02",x"bf",x"6e"),
   265 => (x"74",x"4b",x"87",x"c5"),
   266 => (x"c0",x"0f",x"73",x"49"),
   267 => (x"1e",x"f0",x"c3",x"1e"),
   268 => (x"f6",x"49",x"da",x"c1"),
   269 => (x"86",x"c8",x"87",x"d5"),
   270 => (x"c0",x"02",x"98",x"70"),
   271 => (x"ef",x"c2",x"87",x"d8"),
   272 => (x"6e",x"7e",x"bf",x"c1"),
   273 => (x"c4",x"91",x"cb",x"49"),
   274 => (x"82",x"71",x"4a",x"66"),
   275 => (x"c5",x"c0",x"02",x"6a"),
   276 => (x"49",x"6e",x"4b",x"87"),
   277 => (x"9d",x"75",x"0f",x"73"),
   278 => (x"87",x"c8",x"c0",x"02"),
   279 => (x"bf",x"c1",x"ef",x"c2"),
   280 => (x"87",x"eb",x"f1",x"49"),
   281 => (x"bf",x"fc",x"d3",x"c2"),
   282 => (x"87",x"dd",x"c0",x"02"),
   283 => (x"87",x"dc",x"c2",x"49"),
   284 => (x"c0",x"02",x"98",x"70"),
   285 => (x"ef",x"c2",x"87",x"d3"),
   286 => (x"f1",x"49",x"bf",x"c1"),
   287 => (x"49",x"c0",x"87",x"d1"),
   288 => (x"c2",x"87",x"f1",x"f2"),
   289 => (x"c0",x"48",x"fc",x"d3"),
   290 => (x"f2",x"8e",x"f8",x"78"),
   291 => (x"5e",x"0e",x"87",x"cb"),
   292 => (x"0e",x"5d",x"5c",x"5b"),
   293 => (x"c2",x"4c",x"71",x"1e"),
   294 => (x"49",x"bf",x"fd",x"ee"),
   295 => (x"4d",x"a1",x"cd",x"c1"),
   296 => (x"69",x"81",x"d1",x"c1"),
   297 => (x"02",x"9c",x"74",x"7e"),
   298 => (x"a5",x"c4",x"87",x"cf"),
   299 => (x"c2",x"7b",x"74",x"4b"),
   300 => (x"49",x"bf",x"fd",x"ee"),
   301 => (x"6e",x"87",x"ea",x"f1"),
   302 => (x"05",x"9c",x"74",x"7b"),
   303 => (x"4b",x"c0",x"87",x"c4"),
   304 => (x"4b",x"c1",x"87",x"c2"),
   305 => (x"eb",x"f1",x"49",x"73"),
   306 => (x"02",x"66",x"d4",x"87"),
   307 => (x"c0",x"49",x"87",x"c8"),
   308 => (x"4a",x"70",x"87",x"ee"),
   309 => (x"4a",x"c0",x"87",x"c2"),
   310 => (x"5a",x"c0",x"d4",x"c2"),
   311 => (x"87",x"f9",x"f0",x"26"),
   312 => (x"00",x"00",x"00",x"00"),
   313 => (x"14",x"11",x"12",x"58"),
   314 => (x"23",x"1c",x"1b",x"1d"),
   315 => (x"94",x"91",x"59",x"5a"),
   316 => (x"f4",x"eb",x"f2",x"f5"),
   317 => (x"00",x"00",x"00",x"00"),
   318 => (x"00",x"00",x"00",x"00"),
   319 => (x"00",x"00",x"00",x"00"),
   320 => (x"ff",x"4a",x"71",x"1e"),
   321 => (x"72",x"49",x"bf",x"c8"),
   322 => (x"4f",x"26",x"48",x"a1"),
   323 => (x"bf",x"c8",x"ff",x"1e"),
   324 => (x"c0",x"c0",x"fe",x"89"),
   325 => (x"a9",x"c0",x"c0",x"c0"),
   326 => (x"c0",x"87",x"c4",x"01"),
   327 => (x"c1",x"87",x"c2",x"4a"),
   328 => (x"26",x"48",x"72",x"4a"),
   329 => (x"5b",x"5e",x"0e",x"4f"),
   330 => (x"71",x"0e",x"5d",x"5c"),
   331 => (x"4c",x"d4",x"ff",x"4b"),
   332 => (x"c0",x"48",x"66",x"d0"),
   333 => (x"ff",x"49",x"d6",x"78"),
   334 => (x"c3",x"87",x"fd",x"da"),
   335 => (x"49",x"6c",x"7c",x"ff"),
   336 => (x"71",x"99",x"ff",x"c3"),
   337 => (x"f0",x"c3",x"49",x"4d"),
   338 => (x"a9",x"e0",x"c1",x"99"),
   339 => (x"c3",x"87",x"cb",x"05"),
   340 => (x"48",x"6c",x"7c",x"ff"),
   341 => (x"66",x"d0",x"98",x"c3"),
   342 => (x"ff",x"c3",x"78",x"08"),
   343 => (x"49",x"4a",x"6c",x"7c"),
   344 => (x"ff",x"c3",x"31",x"c8"),
   345 => (x"71",x"4a",x"6c",x"7c"),
   346 => (x"c8",x"49",x"72",x"b2"),
   347 => (x"7c",x"ff",x"c3",x"31"),
   348 => (x"b2",x"71",x"4a",x"6c"),
   349 => (x"31",x"c8",x"49",x"72"),
   350 => (x"6c",x"7c",x"ff",x"c3"),
   351 => (x"ff",x"b2",x"71",x"4a"),
   352 => (x"e0",x"c0",x"48",x"d0"),
   353 => (x"02",x"9b",x"73",x"78"),
   354 => (x"7b",x"72",x"87",x"c2"),
   355 => (x"4d",x"26",x"48",x"75"),
   356 => (x"4b",x"26",x"4c",x"26"),
   357 => (x"26",x"1e",x"4f",x"26"),
   358 => (x"5b",x"5e",x"0e",x"4f"),
   359 => (x"86",x"f8",x"0e",x"5c"),
   360 => (x"a6",x"c8",x"1e",x"76"),
   361 => (x"87",x"fd",x"fd",x"49"),
   362 => (x"4b",x"70",x"86",x"c4"),
   363 => (x"a8",x"c2",x"48",x"6e"),
   364 => (x"87",x"f0",x"c2",x"03"),
   365 => (x"f0",x"c3",x"4a",x"73"),
   366 => (x"aa",x"d0",x"c1",x"9a"),
   367 => (x"c1",x"87",x"c7",x"02"),
   368 => (x"c2",x"05",x"aa",x"e0"),
   369 => (x"49",x"73",x"87",x"de"),
   370 => (x"c3",x"02",x"99",x"c8"),
   371 => (x"87",x"c6",x"ff",x"87"),
   372 => (x"9c",x"c3",x"4c",x"73"),
   373 => (x"c1",x"05",x"ac",x"c2"),
   374 => (x"66",x"c4",x"87",x"c2"),
   375 => (x"71",x"31",x"c9",x"49"),
   376 => (x"4a",x"66",x"c4",x"1e"),
   377 => (x"ef",x"c2",x"92",x"d4"),
   378 => (x"81",x"72",x"49",x"c5"),
   379 => (x"87",x"e1",x"cf",x"fe"),
   380 => (x"d8",x"ff",x"49",x"d8"),
   381 => (x"c0",x"c8",x"87",x"c2"),
   382 => (x"e2",x"dd",x"c2",x"1e"),
   383 => (x"dd",x"eb",x"fd",x"49"),
   384 => (x"48",x"d0",x"ff",x"87"),
   385 => (x"c2",x"78",x"e0",x"c0"),
   386 => (x"cc",x"1e",x"e2",x"dd"),
   387 => (x"92",x"d4",x"4a",x"66"),
   388 => (x"49",x"c5",x"ef",x"c2"),
   389 => (x"cd",x"fe",x"81",x"72"),
   390 => (x"86",x"cc",x"87",x"e8"),
   391 => (x"c1",x"05",x"ac",x"c1"),
   392 => (x"66",x"c4",x"87",x"c2"),
   393 => (x"71",x"31",x"c9",x"49"),
   394 => (x"4a",x"66",x"c4",x"1e"),
   395 => (x"ef",x"c2",x"92",x"d4"),
   396 => (x"81",x"72",x"49",x"c5"),
   397 => (x"87",x"d9",x"ce",x"fe"),
   398 => (x"1e",x"e2",x"dd",x"c2"),
   399 => (x"d4",x"4a",x"66",x"c8"),
   400 => (x"c5",x"ef",x"c2",x"92"),
   401 => (x"fe",x"81",x"72",x"49"),
   402 => (x"d7",x"87",x"e8",x"cb"),
   403 => (x"e7",x"d6",x"ff",x"49"),
   404 => (x"1e",x"c0",x"c8",x"87"),
   405 => (x"49",x"e2",x"dd",x"c2"),
   406 => (x"87",x"db",x"e9",x"fd"),
   407 => (x"d0",x"ff",x"86",x"cc"),
   408 => (x"78",x"e0",x"c0",x"48"),
   409 => (x"e7",x"fc",x"8e",x"f8"),
   410 => (x"5b",x"5e",x"0e",x"87"),
   411 => (x"1e",x"0e",x"5d",x"5c"),
   412 => (x"d4",x"ff",x"4d",x"71"),
   413 => (x"7e",x"66",x"d4",x"4c"),
   414 => (x"a8",x"b7",x"c3",x"48"),
   415 => (x"c0",x"87",x"c5",x"06"),
   416 => (x"87",x"e2",x"c1",x"48"),
   417 => (x"dc",x"fe",x"49",x"75"),
   418 => (x"1e",x"75",x"87",x"d4"),
   419 => (x"d4",x"4b",x"66",x"c4"),
   420 => (x"c5",x"ef",x"c2",x"93"),
   421 => (x"fe",x"49",x"73",x"83"),
   422 => (x"c8",x"87",x"e5",x"c5"),
   423 => (x"ff",x"4b",x"6b",x"83"),
   424 => (x"e1",x"c8",x"48",x"d0"),
   425 => (x"73",x"7c",x"dd",x"78"),
   426 => (x"99",x"ff",x"c3",x"49"),
   427 => (x"49",x"73",x"7c",x"71"),
   428 => (x"c3",x"29",x"b7",x"c8"),
   429 => (x"7c",x"71",x"99",x"ff"),
   430 => (x"b7",x"d0",x"49",x"73"),
   431 => (x"99",x"ff",x"c3",x"29"),
   432 => (x"49",x"73",x"7c",x"71"),
   433 => (x"71",x"29",x"b7",x"d8"),
   434 => (x"7c",x"7c",x"c0",x"7c"),
   435 => (x"7c",x"7c",x"7c",x"7c"),
   436 => (x"7c",x"7c",x"7c",x"7c"),
   437 => (x"e0",x"c0",x"7c",x"7c"),
   438 => (x"1e",x"66",x"c4",x"78"),
   439 => (x"d4",x"ff",x"49",x"dc"),
   440 => (x"86",x"c8",x"87",x"fb"),
   441 => (x"fa",x"26",x"48",x"73"),
   442 => (x"73",x"1e",x"87",x"e4"),
   443 => (x"c2",x"4b",x"c0",x"1e"),
   444 => (x"c0",x"48",x"ef",x"dc"),
   445 => (x"eb",x"dc",x"c2",x"50"),
   446 => (x"de",x"fe",x"49",x"bf"),
   447 => (x"98",x"70",x"87",x"c4"),
   448 => (x"c2",x"87",x"c4",x"05"),
   449 => (x"73",x"4b",x"d3",x"dc"),
   450 => (x"26",x"87",x"c4",x"48"),
   451 => (x"26",x"4c",x"26",x"4d"),
   452 => (x"53",x"4f",x"26",x"4b"),
   453 => (x"2f",x"77",x"6f",x"68"),
   454 => (x"65",x"64",x"69",x"68"),
   455 => (x"44",x"53",x"4f",x"20"),
   456 => (x"6b",x"20",x"3d",x"20"),
   457 => (x"46",x"20",x"79",x"65"),
   458 => (x"30",x"00",x"32",x"31"),
   459 => (x"00",x"00",x"00",x"27"),
   460 => (x"4f",x"54",x"55",x"41"),
   461 => (x"54",x"4f",x"4f",x"42"),
   462 => (x"00",x"53",x"45",x"4e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

